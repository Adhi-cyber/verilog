module t_ff(clk, t, rst, q);

input clk;
input t;
input rst;

output reg q;

always @(posedge clk)
	begin
		if(!rst)
			q <= 0;
		else 
			if(t)
				q <= ~q;
			else
				q <= q;
		end
		endmodule
