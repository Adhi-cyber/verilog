module block_assign_des_2(din, clk, a, b, c);

input din;
input clk;

output reg a;
output reg b;
output reg c;

always @(posedge clk)
begin
        b = a;
        c = b;
	a = din;

end
endmodule

module block_assign_tes_2;

reg din;
reg clk;

wire a;
wire b;
wire c;

block_assign_des_2 uut(.din(din),
        .clk(clk),
        .a(a),
        .b(b),
        .c(c));

initial
begin
        $dumpfile("block_wave_2.vcd");
        $dumpvars(0,block_assign_tes_2);
        din = 1'b1;
        clk = 1'b0;
end

always #2 clk = clk + 1'b1;

endmodule

















































































































































































































































































































































































































































































































































































































































































































































































